/**
* Author: YangHui
* Date: 20220401
* File: clint.v
*/

`ifndef __ISE__
`include "rtl/core/define.v"
`endif

`ifdef __ISE__
`include "define.v"
`endif

module clint (

);
    
endmodule