/**
* Author: YangHui
* Date: 20220401
* File: clint.v
*/

`ifndef __ISE__
`include "rtl/core/define.v"
`endif

module clint (

);
    
endmodule