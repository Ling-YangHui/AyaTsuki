/** 
* Author: YangHui
* Date: 20220403
* File: bus.v
*/

`ifndef __ISE__
`include "rtl/core/define.v"
`endif

module bus (
    
);
    
endmodule